`timescale 1ns/1ns
module Shifter( dataA, dataB, Signal, dataOut, reset );
input reset ;
input [31:0] dataA ;
input [4:0] dataB ;     // 移位量
input [5:0] Signal ;
output [31:0] dataOut ;
wire [31:0] s0,s1,s2,s3,s4 ; // 每層之間的接線 
wire [31:0] temp ;

parameter SLL = 6'b000000;
    
  // 左移一位元
  mux2to1 m1_0 ( 1'b0    , dataA[0], s0[0], dataB[0] ) ;
  mux2to1 m1_1 ( dataA[0], dataA[1], s0[1], dataB[0] ) ;
  mux2to1 m1_2 ( dataA[1], dataA[2], s0[2], dataB[0] ) ;
  mux2to1 m1_3 ( dataA[2], dataA[3], s0[3], dataB[0] ) ;
  mux2to1 m1_4 ( dataA[3], dataA[4], s0[4], dataB[0] ) ;
  mux2to1 m1_5 ( dataA[4], dataA[5], s0[5], dataB[0] ) ;
  mux2to1 m1_6 ( dataA[5], dataA[6], s0[6], dataB[0] ) ;
  mux2to1 m1_7 ( dataA[6], dataA[7], s0[7], dataB[0] ) ;
  mux2to1 m1_8 ( dataA[7], dataA[8], s0[8], dataB[0] ) ;
  mux2to1 m1_9 ( dataA[8], dataA[9], s0[9], dataB[0] ) ;
  mux2to1 m1_10 ( dataA[9] , dataA[10], s0[10], dataB[0] ) ;
  mux2to1 m1_11 ( dataA[10], dataA[11], s0[11], dataB[0] ) ;
  mux2to1 m1_12 ( dataA[11], dataA[12], s0[12], dataB[0] ) ;
  mux2to1 m1_13 ( dataA[12], dataA[13], s0[13], dataB[0] ) ;
  mux2to1 m1_14 ( dataA[13], dataA[14], s0[14], dataB[0] ) ;
  mux2to1 m1_15 ( dataA[14], dataA[15], s0[15], dataB[0] ) ;
  mux2to1 m1_16 ( dataA[15], dataA[16], s0[16], dataB[0] ) ;
  mux2to1 m1_17 ( dataA[16], dataA[17], s0[17], dataB[0] ) ;
  mux2to1 m1_18 ( dataA[17], dataA[18], s0[18], dataB[0] ) ;
  mux2to1 m1_19 ( dataA[18], dataA[19], s0[19], dataB[0] ) ;
  mux2to1 m1_20 ( dataA[19], dataA[20], s0[20], dataB[0] ) ;
  mux2to1 m1_21 ( dataA[20], dataA[21], s0[21], dataB[0] ) ;
  mux2to1 m1_22 ( dataA[21], dataA[22], s0[22], dataB[0] ) ;
  mux2to1 m1_23 ( dataA[22], dataA[23], s0[23], dataB[0] ) ;
  mux2to1 m1_24 ( dataA[23], dataA[24], s0[24], dataB[0] ) ;
  mux2to1 m1_25 ( dataA[24], dataA[25], s0[25], dataB[0] ) ;
  mux2to1 m1_26 ( dataA[25], dataA[26], s0[26], dataB[0] ) ;
  mux2to1 m1_27 ( dataA[26], dataA[27], s0[27], dataB[0] ) ;
  mux2to1 m1_28 ( dataA[27], dataA[28], s0[28], dataB[0] ) ;
  mux2to1 m1_29 ( dataA[28], dataA[29], s0[29], dataB[0] ) ;
  mux2to1 m1_30 ( dataA[29], dataA[30], s0[30], dataB[0] ) ;
  mux2to1 m1_31 ( dataA[30], dataA[31], s0[31], dataB[0] ) ;
  // 左移二位元
  mux2to1 m2_0 ( 1'b0, s0[0], s1[0], dataB[1] ) ;
  mux2to1 m2_1 ( 1'b0, s0[1], s1[1], dataB[1] ) ;
  mux2to1 m2_2 ( s0[0], s0[2], s1[2], dataB[1] ) ;
  mux2to1 m2_3 ( s0[1], s0[3], s1[3], dataB[1] ) ;
  mux2to1 m2_4 ( s0[2], s0[4], s1[4], dataB[1] ) ;
  mux2to1 m2_5 ( s0[3], s0[5], s1[5], dataB[1] ) ;
  mux2to1 m2_6 ( s0[4], s0[6], s1[6], dataB[1] ) ;
  mux2to1 m2_7 ( s0[5], s0[7], s1[7], dataB[1] ) ;
  mux2to1 m2_8 ( s0[6], s0[8], s1[8], dataB[1] ) ;
  mux2to1 m2_9 ( s0[7], s0[9], s1[9], dataB[1] ) ;
  mux2to1 m2_10 ( s0[8], s0[10], s1[10], dataB[1] ) ;
  mux2to1 m2_11 ( s0[9], s0[11], s1[11], dataB[1] ) ;
  mux2to1 m2_12 ( s0[10], s0[12], s1[12], dataB[1] ) ;
  mux2to1 m2_13 ( s0[11], s0[13], s1[13], dataB[1] ) ;
  mux2to1 m2_14 ( s0[12], s0[14], s1[14], dataB[1] ) ;
  mux2to1 m2_15 ( s0[13], s0[15], s1[15], dataB[1] ) ;
  mux2to1 m2_16 ( s0[14], s0[16], s1[16], dataB[1] ) ;
  mux2to1 m2_17 ( s0[15], s0[17], s1[17], dataB[1] ) ;
  mux2to1 m2_18 ( s0[16], s0[18], s1[18], dataB[1] ) ;
  mux2to1 m2_19 ( s0[17], s0[19], s1[19], dataB[1] ) ;
  mux2to1 m2_20 ( s0[18], s0[20], s1[20], dataB[1] ) ;
  mux2to1 m2_21 ( s0[19], s0[21], s1[21], dataB[1] ) ;
  mux2to1 m2_22 ( s0[20], s0[22], s1[22], dataB[1] ) ;
  mux2to1 m2_23 ( s0[21], s0[23], s1[23], dataB[1] ) ;
  mux2to1 m2_24 ( s0[22], s0[24], s1[24], dataB[1] ) ;
  mux2to1 m2_25 ( s0[23], s0[25], s1[25], dataB[1] ) ;
  mux2to1 m2_26 ( s0[24], s0[26], s1[26], dataB[1] ) ;
  mux2to1 m2_27 ( s0[25], s0[27], s1[27], dataB[1] ) ;
  mux2to1 m2_28 ( s0[26], s0[28], s1[28], dataB[1] ) ;
  mux2to1 m2_29 ( s0[27], s0[29], s1[29], dataB[1] ) ;
  mux2to1 m2_30 ( s0[28], s0[30], s1[30], dataB[1] ) ;
  mux2to1 m2_31 ( s0[29], s0[31], s1[31], dataB[1] ) ;
  // 左移四位元
  mux2to1 m3_0 ( 1'b0, s1[0], s2[0], dataB[2] ) ;
  mux2to1 m3_1 ( 1'b0, s1[1], s2[1], dataB[2] ) ;
  mux2to1 m3_2 ( 1'b0, s1[2], s2[2], dataB[2] ) ;
  mux2to1 m3_3 ( 1'b0, s1[3], s2[3], dataB[2] ) ;
  mux2to1 m3_4 ( s1[0], s1[4], s2[4], dataB[2] ) ;
  mux2to1 m3_5 ( s1[1], s1[5], s2[5], dataB[2] ) ;
  mux2to1 m3_6 ( s1[2], s1[6], s2[6], dataB[2] ) ;
  mux2to1 m3_7 ( s1[3], s1[7], s2[7], dataB[2] ) ;
  mux2to1 m3_8 ( s1[4], s1[8], s2[8], dataB[2] ) ;
  mux2to1 m3_9 ( s1[5], s1[9], s2[9], dataB[2] ) ;
  mux2to1 m3_10 ( s1[6], s1[10], s2[10], dataB[2] ) ;
  mux2to1 m3_11 ( s1[7], s1[11], s2[11], dataB[2] ) ;
  mux2to1 m3_12 ( s1[8], s1[12], s2[12], dataB[2] ) ;
  mux2to1 m3_13 ( s1[9], s1[13], s2[13], dataB[2] ) ;
  mux2to1 m3_14 ( s1[10], s1[14], s2[14], dataB[2] ) ;
  mux2to1 m3_15 ( s1[11], s1[15], s2[15], dataB[2] ) ;
  mux2to1 m3_16 ( s1[12], s1[16], s2[16], dataB[2] ) ;
  mux2to1 m3_17 ( s1[13], s1[17], s2[17], dataB[2] ) ;
  mux2to1 m3_18 ( s1[14], s1[18], s2[18], dataB[2] ) ;
  mux2to1 m3_19 ( s1[15], s1[19], s2[19], dataB[2] ) ;
  mux2to1 m3_20 ( s1[16], s1[20], s2[20], dataB[2] ) ;
  mux2to1 m3_21 ( s1[17], s1[21], s2[21], dataB[2] ) ;
  mux2to1 m3_22 ( s1[18], s1[22], s2[22], dataB[2] ) ;
  mux2to1 m3_23 ( s1[19], s1[23], s2[23], dataB[2] ) ;
  mux2to1 m3_24 ( s1[20], s1[24], s2[24], dataB[2] ) ;
  mux2to1 m3_25 ( s1[21], s1[25], s2[25], dataB[2] ) ;
  mux2to1 m3_26 ( s1[22], s1[26], s2[26], dataB[2] ) ;
  mux2to1 m3_27 ( s1[23], s1[27], s2[27], dataB[2] ) ;
  mux2to1 m3_28 ( s1[24], s1[28], s2[28], dataB[2] ) ;
  mux2to1 m3_29 ( s1[25], s1[29], s2[29], dataB[2] ) ;
  mux2to1 m3_30 ( s1[26], s1[30], s2[30], dataB[2] ) ;
  mux2to1 m3_31 ( s1[27], s1[31], s2[31], dataB[2] ) ;
  // 左移八位元
  mux2to1 m4_0 ( 1'b0, s2[0], s3[0], dataB[3] ) ;
  mux2to1 m4_1 ( 1'b0, s2[1], s3[1], dataB[3] ) ;
  mux2to1 m4_2 ( 1'b0, s2[2], s3[2], dataB[3] ) ;
  mux2to1 m4_3 ( 1'b0, s2[3], s3[3], dataB[3] ) ;
  mux2to1 m4_4 ( 1'b0, s2[4], s3[4], dataB[3] ) ;
  mux2to1 m4_5 ( 1'b0, s2[5], s3[5], dataB[3] ) ;
  mux2to1 m4_6 ( 1'b0, s2[6], s3[6], dataB[3] ) ;
  mux2to1 m4_7 ( 1'b0, s2[7], s3[7], dataB[3] ) ;
  mux2to1 m4_8 ( s2[0], s2[8], s3[8], dataB[3] ) ;
  mux2to1 m4_9 ( s2[1], s2[9], s3[9], dataB[3] ) ;
  mux2to1 m4_10 ( s2[2], s2[10], s3[10], dataB[3] ) ;
  mux2to1 m4_11 ( s2[3], s2[11], s3[11], dataB[3] ) ;
  mux2to1 m4_12 ( s2[4], s2[12], s3[12], dataB[3] ) ;
  mux2to1 m4_13 ( s2[5], s2[13], s3[13], dataB[3] ) ;
  mux2to1 m4_14 ( s2[6], s2[14], s3[14], dataB[3] ) ;
  mux2to1 m4_15 ( s2[7], s2[15], s3[15], dataB[3] ) ;
  mux2to1 m4_16 ( s2[8], s2[16], s3[16], dataB[3] ) ;
  mux2to1 m4_17 ( s2[9], s2[17], s3[17], dataB[3] ) ;
  mux2to1 m4_18 ( s2[10], s2[18], s3[18], dataB[3] ) ;
  mux2to1 m4_19 ( s2[11], s2[19], s3[19], dataB[3] ) ;
  mux2to1 m4_20 ( s2[12], s2[20], s3[20], dataB[3] ) ;
  mux2to1 m4_21 ( s2[13], s2[21], s3[21], dataB[3] ) ;
  mux2to1 m4_22 ( s2[14], s2[22], s3[22], dataB[3] ) ;
  mux2to1 m4_23 ( s2[15], s2[23], s3[23], dataB[3] ) ;
  mux2to1 m4_24 ( s2[16], s2[24], s3[24], dataB[3] ) ;
  mux2to1 m4_25 ( s2[17], s2[25], s3[25], dataB[3] ) ;
  mux2to1 m4_26 ( s2[18], s2[26], s3[26], dataB[3] ) ;
  mux2to1 m4_27 ( s2[19], s2[27], s3[27], dataB[3] ) ;
  mux2to1 m4_28 ( s2[20], s2[28], s3[28], dataB[3] ) ;
  mux2to1 m4_29 ( s2[21], s2[29], s3[29], dataB[3] ) ;
  mux2to1 m4_30 ( s2[22], s2[30], s3[30], dataB[3] ) ;
  mux2to1 m4_31 ( s2[23], s2[31], s3[31], dataB[3] ) ;
  // 左移16位元
  mux2to1 m5_0 ( 1'b0, s3[0], s4[0], dataB[4] ) ;
  mux2to1 m5_1 ( 1'b0, s3[1], s4[1], dataB[4] ) ;
  mux2to1 m5_2 ( 1'b0, s3[2], s4[2], dataB[4] ) ;
  mux2to1 m5_3 ( 1'b0, s3[3], s4[3], dataB[4] ) ;
  mux2to1 m5_4 ( 1'b0, s3[4], s4[4], dataB[4] ) ;
  mux2to1 m5_5 ( 1'b0, s3[5], s4[5], dataB[4] ) ;
  mux2to1 m5_6 ( 1'b0, s3[6], s4[6], dataB[4] ) ;
  mux2to1 m5_7 ( 1'b0, s3[7], s4[7], dataB[4] ) ;
  mux2to1 m5_8 ( 1'b0, s3[8], s4[8], dataB[4] ) ;
  mux2to1 m5_9 ( 1'b0, s3[9], s4[9], dataB[4] ) ;
  mux2to1 m5_10 ( 1'b0, s3[10], s4[10], dataB[4] ) ;
  mux2to1 m5_11 ( 1'b0, s3[11], s4[11], dataB[4] ) ;
  mux2to1 m5_12 ( 1'b0, s3[12], s4[12], dataB[4] ) ;
  mux2to1 m5_13 ( 1'b0, s3[13], s4[13], dataB[4] ) ;
  mux2to1 m5_14 ( 1'b0, s3[14], s4[14], dataB[4] ) ;
  mux2to1 m5_15 ( 1'b0, s3[15], s4[15], dataB[4] ) ;
  mux2to1 m5_16 ( s3[0], s3[16], s4[16], dataB[4] ) ;
  mux2to1 m5_17 ( s3[1], s3[17], s4[17], dataB[4] ) ;
  mux2to1 m5_18 ( s3[2], s3[18], s4[18], dataB[4] ) ;
  mux2to1 m5_19 ( s3[3], s3[19], s4[19], dataB[4] ) ;
  mux2to1 m5_20 ( s3[4], s3[20], s4[20], dataB[4] ) ;
  mux2to1 m5_21 ( s3[5], s3[21], s4[21], dataB[4] ) ;
  mux2to1 m5_22 ( s3[6], s3[22], s4[22], dataB[4] ) ;
  mux2to1 m5_23 ( s3[7], s3[23], s4[23], dataB[4] ) ;
  mux2to1 m5_24 ( s3[8], s3[24], s4[24], dataB[4] ) ;
  mux2to1 m5_25 ( s3[9], s3[25], s4[25], dataB[4] ) ;
  mux2to1 m5_26 ( s3[10], s3[26], s4[26], dataB[4] ) ;
  mux2to1 m5_27 ( s3[11], s3[27], s4[27], dataB[4] ) ;
  mux2to1 m5_28 ( s3[12], s3[28], s4[28], dataB[4] ) ;
  mux2to1 m5_29 ( s3[13], s3[29], s4[29], dataB[4] ) ;
  mux2to1 m5_30 ( s3[14], s3[30], s4[30], dataB[4] ) ;
  mux2to1 m5_31 ( s3[15], s3[31], s4[31], dataB[4] ) ;
  
  //  assign temp = ( dataB < 5'd32 ) ? s4 : 0 ;
  assign temp =  s4 ;
  assign dataOut = ( reset ) ? 0 : temp ;
  
endmodule  
  